module mux32_2_1(R, S, A, B);

output [31:0] R;
input S;
input [31:0] A, B;

	mux_2_1 m31(R[31], S, A[31], B[31]);
	mux_2_1 m30(R[30], S, A[30], B[30]);
	mux_2_1 m29(R[29], S, A[29], B[29]);
	mux_2_1 m28(R[28], S, A[28], B[28]);
	mux_2_1 m27(R[27], S, A[27], B[27]);
	mux_2_1 m26(R[26], S, A[26], B[26]);
	mux_2_1 m25(R[25], S, A[25], B[25]);
	mux_2_1 m24(R[24], S, A[24], B[24]);
	mux_2_1 m23(R[23], S, A[23], B[23]);
	mux_2_1 m22(R[22], S, A[22], B[22]);
	mux_2_1 m21(R[21], S, A[21], B[21]);
	mux_2_1 m20(R[20], S, A[20], B[20]);
	mux_2_1 m19(R[19], S, A[19], B[19]);
	mux_2_1 m18(R[18], S, A[18], B[18]);
	mux_2_1 m17(R[17], S, A[17], B[17]);
	mux_2_1 m16(R[16], S, A[16], B[16]);
	mux_2_1 m15(R[15], S, A[15], B[15]);
	mux_2_1 m14(R[14], S, A[14], B[14]);
	mux_2_1 m13(R[13], S, A[13], B[13]);
	mux_2_1 m12(R[12], S, A[12], B[12]);
	mux_2_1 m11(R[11], S, A[11], B[11]);
	mux_2_1 m10(R[10], S, A[10], B[10]);
	mux_2_1 m9 (R[9],  S, A[9],  B[9]);
	mux_2_1 m8 (R[8],  S, A[8],  B[8]);
	mux_2_1 m7 (R[7],  S, A[7],  B[7]);
	mux_2_1 m6 (R[6],  S, A[6],  B[6]);
	mux_2_1 m5 (R[5],  S, A[5],  B[5]);
	mux_2_1 m4 (R[4],  S, A[4],  B[4]);
	mux_2_1 m3 (R[3],  S, A[3],  B[3]);
	mux_2_1 m2 (R[2],  S, A[2],  B[2]);
	mux_2_1 m1 (R[1],  S, A[1],  B[1]);
	mux_2_1 m0 (R[0],  S, A[0],  B[0]);
	

endmodule 
