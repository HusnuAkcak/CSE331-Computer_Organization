`timescale 1 ps / 1 ps
module sub_32_tb();

	reg [31:0] A, B;
	wire [31:0] R;

	reg clk;

	sub_32 sub_32_inst(R, A, B);
	
	always
		begin 
			#1 clk = ~clk;
		end
		
	initial 
		begin 
			A = 32'b00000000000000000000000000000111; //7
			B = 32'b00000000000000000000000000100000; //32
			// 7-32 => 25 => 32'b11111111111111111111111111100111
			
		 #100 
			A = 32'b00000000000000000000000000001111; //15
			B = 32'b00000000000000000000000000010000; //16
			// 15-16 => 17 => 32'b11111111111111111111111111111111
	
		#100 
			A = 32'b00000000000000000000000000000101; // 5
			B = 32'b11111111111111111111111111111101;	// -3		 
			// 5-(-3) => 8 => 32'b00000000000000000000000000001000

		#100 
			A = 32'b00000000000000000000000000000101; //5
			B = 32'b00000000000000000000000000000100; //4
			// 5-4 => 1 => 32'b00000000000000000000000000000001
			
			
		end
		
		initial begin
		$monitor("time = %2d\n A = %32b\n B = %32b\n R = %32b \n\n",
				$time, A, B, R);
		end
	
endmodule
