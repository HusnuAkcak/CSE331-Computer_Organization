`timescale 1 ps / 1 ps
module slt_32_tb();

	reg [31:0] A, B;
	wire [31:0] R;

	reg clk;

	slt_32 slt_32_inst(R, A, B);
	
	always
		begin 
			#1 clk = ~clk;
		end
		
	initial 
		begin 
			A = 32'b00000000000000000000000000000111; // 7
			B = 32'b00000000000000000000000000100000; // 32
			
		 #100 
			A = 32'b00000000000000000000000000001111; // 15
			B = 32'b00000000000000000000000000010000; // 16
	
		#100 
			A = 32'b00000000000000000000000000000101; // 5
			B = 32'b11111111111111111111111111111101;	// -3		 

		#100 
			A = 32'b00000000000000000000000000000101; // 5
			B = 32'b00000000000000000000000000000100; // 4
			
		
		#100 
			A = 32'b11111111111111111111111111111100; // -4
			B = 32'b11111111111111111111111111111101;	// -3		 

			
		#100 
			A = 32'b11111111111111111111111111111101;	// -3		
			B = 32'b11111111111111111111111111111100; // -4 

			
		end
		
		initial begin
		$monitor("time = %2d\n A = %32b\n B = %32b\n R = %32b \n\n",
				$time, A, B, R);
		end
	
endmodule
